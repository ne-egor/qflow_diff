VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 1.900 0.000 ;
  SIZE 66.200 BY 44.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.400 40.400 57.200 41.600 ;
        RECT 2.800 33.000 3.600 40.400 ;
        RECT 6.000 31.800 6.800 40.400 ;
        RECT 15.600 35.800 16.400 40.400 ;
        RECT 18.800 32.200 19.600 40.400 ;
        RECT 22.000 35.800 22.800 40.400 ;
        RECT 25.200 35.800 26.000 40.400 ;
        RECT 28.400 35.800 29.200 40.400 ;
        RECT 31.600 35.800 32.400 40.400 ;
        RECT 39.600 35.800 40.400 40.400 ;
        RECT 42.800 35.800 43.600 40.400 ;
        RECT 49.200 35.800 50.000 40.400 ;
        RECT 52.400 35.800 53.200 40.400 ;
        RECT 55.600 35.800 56.400 40.400 ;
        RECT 49.000 31.800 49.800 32.000 ;
        RECT 52.400 31.800 53.200 32.400 ;
        RECT 26.200 31.200 53.200 31.800 ;
        RECT 26.200 31.000 27.000 31.200 ;
        RECT 23.000 10.800 23.800 11.000 ;
        RECT 23.000 10.200 50.000 10.800 ;
        RECT 2.800 1.600 3.600 9.000 ;
        RECT 6.000 1.600 6.800 6.200 ;
        RECT 9.200 1.600 10.000 10.200 ;
        RECT 45.800 10.000 46.600 10.200 ;
        RECT 49.200 9.600 50.000 10.200 ;
        RECT 18.800 1.600 19.600 6.200 ;
        RECT 22.000 1.600 22.800 6.200 ;
        RECT 25.200 1.600 26.000 6.200 ;
        RECT 28.400 1.600 29.200 6.200 ;
        RECT 36.400 1.600 37.200 6.200 ;
        RECT 39.600 1.600 40.400 6.200 ;
        RECT 46.000 1.600 46.800 6.200 ;
        RECT 49.200 1.600 50.000 6.200 ;
        RECT 52.400 1.600 53.200 6.200 ;
        RECT 60.400 1.600 61.200 6.200 ;
        RECT 0.400 0.400 62.000 1.600 ;
      LAYER via1 ;
        RECT 12.600 40.600 13.400 41.400 ;
        RECT 14.000 40.600 14.800 41.400 ;
        RECT 15.400 40.600 16.200 41.400 ;
        RECT 52.400 37.600 53.200 38.400 ;
        RECT 52.400 31.600 53.200 32.400 ;
        RECT 49.200 3.600 50.000 4.400 ;
        RECT 12.600 0.600 13.400 1.400 ;
        RECT 14.000 0.600 14.800 1.400 ;
        RECT 15.400 0.600 16.200 1.400 ;
      LAYER metal2 ;
        RECT 12.000 40.600 16.800 41.400 ;
        RECT 52.400 37.600 53.200 38.400 ;
        RECT 52.500 32.400 53.100 37.600 ;
        RECT 52.400 31.600 53.200 32.400 ;
        RECT 49.200 9.600 50.000 10.400 ;
        RECT 49.300 4.400 49.900 9.600 ;
        RECT 49.200 3.600 50.000 4.400 ;
        RECT 12.000 0.600 16.800 1.400 ;
      LAYER via2 ;
        RECT 12.600 40.600 13.400 41.400 ;
        RECT 14.000 40.600 14.800 41.400 ;
        RECT 15.400 40.600 16.200 41.400 ;
        RECT 12.600 0.600 13.400 1.400 ;
        RECT 14.000 0.600 14.800 1.400 ;
        RECT 15.400 0.600 16.200 1.400 ;
      LAYER metal3 ;
        RECT 12.000 40.400 16.800 41.600 ;
        RECT 12.000 0.400 16.800 1.600 ;
      LAYER via3 ;
        RECT 12.400 40.600 13.200 41.400 ;
        RECT 14.000 40.600 14.800 41.400 ;
        RECT 15.600 40.600 16.400 41.400 ;
        RECT 12.400 0.600 13.200 1.400 ;
        RECT 14.000 0.600 14.800 1.400 ;
        RECT 15.600 0.600 16.400 1.400 ;
      LAYER metal4 ;
        RECT 12.000 0.000 16.800 44.000 ;
    END
  END vdd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 38.800 25.600 40.400 26.400 ;
        RECT 35.600 15.600 37.200 16.400 ;
      LAYER via1 ;
        RECT 39.600 25.600 40.400 26.400 ;
        RECT 36.400 15.600 37.200 16.400 ;
      LAYER metal2 ;
        RECT 42.900 40.400 43.500 44.300 ;
        RECT 39.600 39.600 40.400 40.400 ;
        RECT 42.800 39.600 43.600 40.400 ;
        RECT 39.700 26.400 40.300 39.600 ;
        RECT 39.600 25.600 40.400 26.400 ;
        RECT 39.700 16.400 40.300 25.600 ;
        RECT 36.400 15.600 37.200 16.400 ;
        RECT 39.600 15.600 40.400 16.400 ;
      LAYER metal3 ;
        RECT 39.600 40.300 40.400 40.400 ;
        RECT 42.800 40.300 43.600 40.400 ;
        RECT 39.600 39.700 43.600 40.300 ;
        RECT 39.600 39.600 40.400 39.700 ;
        RECT 42.800 39.600 43.600 39.700 ;
        RECT 36.400 16.300 37.200 16.400 ;
        RECT 39.600 16.300 40.400 16.400 ;
        RECT 36.400 15.700 40.400 16.300 ;
        RECT 36.400 15.600 37.200 15.700 ;
        RECT 39.600 15.600 40.400 15.700 ;
    END
  END clk
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 60.400 15.600 61.200 17.200 ;
      LAYER metal2 ;
        RECT 60.400 15.600 61.200 16.400 ;
        RECT 60.500 10.400 61.100 15.600 ;
        RECT 60.400 9.600 61.200 10.400 ;
      LAYER metal3 ;
        RECT 60.400 10.300 61.200 10.400 ;
        RECT 60.400 9.700 64.300 10.300 ;
        RECT 60.400 9.600 61.200 9.700 ;
    END
  END rst
  PIN val[0]
    PORT
      LAYER metal1 ;
        RECT 1.200 12.400 2.000 19.800 ;
        RECT 1.200 10.200 1.800 12.400 ;
        RECT 1.200 2.200 2.000 10.200 ;
      LAYER via1 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal2 ;
        RECT 1.200 9.600 2.000 10.400 ;
        RECT 1.300 8.400 1.900 9.600 ;
        RECT 1.200 7.600 2.000 8.400 ;
      LAYER metal3 ;
        RECT 1.200 10.300 2.000 10.400 ;
        RECT -1.900 9.700 2.000 10.300 ;
        RECT 1.200 9.600 2.000 9.700 ;
    END
  END val[0]
  PIN val[1]
    PORT
      LAYER metal1 ;
        RECT 1.200 31.800 2.000 39.800 ;
        RECT 1.200 29.600 1.800 31.800 ;
        RECT 1.200 22.200 2.000 29.600 ;
      LAYER via1 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal2 ;
        RECT 1.200 29.600 2.000 30.400 ;
        RECT 1.300 28.400 1.900 29.600 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal3 ;
        RECT 1.200 30.300 2.000 30.400 ;
        RECT -1.900 29.700 2.000 30.300 ;
        RECT 1.200 29.600 2.000 29.700 ;
    END
  END val[1]
  OBS
      LAYER metal1 ;
        RECT 4.400 32.400 5.200 39.800 ;
        RECT 8.600 32.600 9.400 39.800 ;
        RECT 17.200 35.800 18.000 39.800 ;
        RECT 3.000 31.800 5.200 32.400 ;
        RECT 7.600 31.800 9.400 32.600 ;
        RECT 3.000 31.200 3.600 31.800 ;
        RECT 2.400 30.400 3.600 31.200 ;
        RECT 3.000 27.400 3.600 30.400 ;
        RECT 4.400 30.300 5.200 30.400 ;
        RECT 6.000 30.300 6.800 30.400 ;
        RECT 4.400 29.700 6.800 30.300 ;
        RECT 4.400 28.800 5.200 29.700 ;
        RECT 6.000 29.600 6.800 29.700 ;
        RECT 7.800 28.400 8.400 31.800 ;
        RECT 17.400 31.600 18.000 35.800 ;
        RECT 20.400 31.800 21.200 39.800 ;
        RECT 23.600 32.000 24.400 39.800 ;
        RECT 26.800 35.200 27.600 39.800 ;
        RECT 9.200 29.600 10.000 31.200 ;
        RECT 17.400 31.000 19.800 31.600 ;
        RECT 17.200 29.600 18.000 30.400 ;
        RECT 7.600 27.600 8.400 28.400 ;
        RECT 15.600 27.600 16.400 29.200 ;
        RECT 17.400 28.800 18.000 29.600 ;
        RECT 17.400 28.200 18.400 28.800 ;
        RECT 17.600 28.000 18.400 28.200 ;
        RECT 19.200 27.600 19.800 31.000 ;
        RECT 20.600 30.400 21.200 31.800 ;
        RECT 20.400 29.600 21.200 30.400 ;
        RECT 3.000 26.800 5.200 27.400 ;
        RECT 2.800 21.600 3.600 26.200 ;
        RECT 4.400 22.200 5.200 26.800 ;
        RECT 6.000 24.800 6.800 26.400 ;
        RECT 7.800 26.300 8.400 27.600 ;
        RECT 19.200 27.400 20.000 27.600 ;
        RECT 17.000 27.000 20.000 27.400 ;
        RECT 15.800 26.800 20.000 27.000 ;
        RECT 15.800 26.400 17.600 26.800 ;
        RECT 9.200 26.300 10.000 26.400 ;
        RECT 7.700 25.700 10.000 26.300 ;
        RECT 15.800 26.200 16.400 26.400 ;
        RECT 20.600 26.200 21.200 29.600 ;
        RECT 7.800 24.200 8.400 25.700 ;
        RECT 9.200 25.600 10.000 25.700 ;
        RECT 6.000 21.600 6.800 24.200 ;
        RECT 7.600 22.200 8.400 24.200 ;
        RECT 9.200 21.600 10.000 24.200 ;
        RECT 15.600 22.200 16.400 26.200 ;
        RECT 18.200 21.600 19.000 26.000 ;
        RECT 19.800 25.200 21.200 26.200 ;
        RECT 23.400 31.200 24.400 32.000 ;
        RECT 25.000 34.600 27.600 35.200 ;
        RECT 25.000 33.000 25.600 34.600 ;
        RECT 30.000 34.400 30.800 39.800 ;
        RECT 33.200 37.000 34.000 39.800 ;
        RECT 34.800 37.000 35.600 39.800 ;
        RECT 36.400 37.000 37.200 39.800 ;
        RECT 31.400 34.400 35.600 35.200 ;
        RECT 28.200 33.600 30.800 34.400 ;
        RECT 38.000 33.600 38.800 39.800 ;
        RECT 41.200 35.000 42.000 39.800 ;
        RECT 44.400 35.000 45.200 39.800 ;
        RECT 46.000 37.000 46.800 39.800 ;
        RECT 47.600 37.000 48.400 39.800 ;
        RECT 50.800 35.200 51.600 39.800 ;
        RECT 54.000 36.400 54.800 39.800 ;
        RECT 54.000 35.800 55.000 36.400 ;
        RECT 54.400 35.200 55.000 35.800 ;
        RECT 49.600 34.400 53.800 35.200 ;
        RECT 54.400 34.600 56.400 35.200 ;
        RECT 41.200 33.600 43.800 34.400 ;
        RECT 44.400 33.800 50.200 34.400 ;
        RECT 53.200 34.000 53.800 34.400 ;
        RECT 33.200 33.000 34.000 33.200 ;
        RECT 25.000 32.400 34.000 33.000 ;
        RECT 36.400 33.000 37.200 33.200 ;
        RECT 44.400 33.000 45.000 33.800 ;
        RECT 50.800 33.200 52.200 33.800 ;
        RECT 53.200 33.200 54.800 34.000 ;
        RECT 36.400 32.400 45.000 33.000 ;
        RECT 46.000 33.000 52.200 33.200 ;
        RECT 46.000 32.600 51.400 33.000 ;
        RECT 46.000 32.400 46.800 32.600 ;
        RECT 23.400 26.800 24.200 31.200 ;
        RECT 25.000 30.600 25.600 32.400 ;
        RECT 24.800 30.000 25.600 30.600 ;
        RECT 31.600 30.000 55.000 30.600 ;
        RECT 24.800 28.000 25.400 30.000 ;
        RECT 31.600 29.400 32.400 30.000 ;
        RECT 49.200 29.600 50.000 30.000 ;
        RECT 54.000 29.800 55.000 30.000 ;
        RECT 54.000 29.600 54.800 29.800 ;
        RECT 26.000 28.600 29.800 29.400 ;
        RECT 24.800 27.400 26.000 28.000 ;
        RECT 23.400 26.000 24.400 26.800 ;
        RECT 19.800 24.400 20.600 25.200 ;
        RECT 19.800 23.600 21.200 24.400 ;
        RECT 19.800 22.200 20.600 23.600 ;
        RECT 22.000 21.600 22.800 24.200 ;
        RECT 23.600 22.200 24.400 26.000 ;
        RECT 25.200 22.200 26.000 27.400 ;
        RECT 29.000 27.400 29.800 28.600 ;
        RECT 29.000 26.800 30.800 27.400 ;
        RECT 30.000 26.200 30.800 26.800 ;
        RECT 34.800 26.400 35.600 29.200 ;
        RECT 38.000 28.600 41.200 29.400 ;
        RECT 45.000 28.600 47.000 29.400 ;
        RECT 55.600 29.000 56.400 34.600 ;
        RECT 37.600 27.800 38.400 28.000 ;
        RECT 37.600 27.200 42.000 27.800 ;
        RECT 41.200 27.000 42.000 27.200 ;
        RECT 42.800 26.800 43.600 28.400 ;
        RECT 28.400 21.600 29.200 26.200 ;
        RECT 30.000 25.400 32.400 26.200 ;
        RECT 34.800 25.600 35.800 26.400 ;
        RECT 41.200 26.200 42.000 26.400 ;
        RECT 45.000 26.200 45.800 28.600 ;
        RECT 47.600 28.200 56.400 29.000 ;
        RECT 51.000 26.800 54.000 27.600 ;
        RECT 51.000 26.200 51.800 26.800 ;
        RECT 41.200 25.600 45.800 26.200 ;
        RECT 31.600 22.200 32.400 25.400 ;
        RECT 49.200 25.400 51.800 26.200 ;
        RECT 33.200 22.200 34.000 25.000 ;
        RECT 34.800 22.200 35.600 25.000 ;
        RECT 36.400 22.200 37.200 25.000 ;
        RECT 38.000 22.200 38.800 25.000 ;
        RECT 39.600 21.600 40.400 24.200 ;
        RECT 41.200 22.200 42.000 25.000 ;
        RECT 42.800 21.600 43.600 24.200 ;
        RECT 44.400 22.200 45.200 25.000 ;
        RECT 46.000 22.200 46.800 25.000 ;
        RECT 47.600 22.200 48.400 25.000 ;
        RECT 49.200 22.200 50.000 25.400 ;
        RECT 52.400 21.600 53.200 26.200 ;
        RECT 55.600 22.200 56.400 28.200 ;
        RECT 0.400 20.400 62.000 21.600 ;
        RECT 2.800 15.800 3.600 20.400 ;
        RECT 4.400 15.200 5.200 19.800 ;
        RECT 6.000 17.800 6.800 20.400 ;
        RECT 6.000 15.600 6.800 17.200 ;
        RECT 3.000 14.600 5.200 15.200 ;
        RECT 3.000 11.600 3.600 14.600 ;
        RECT 4.400 12.300 5.200 13.200 ;
        RECT 6.000 12.300 6.800 12.400 ;
        RECT 4.400 11.700 6.800 12.300 ;
        RECT 4.400 11.600 5.200 11.700 ;
        RECT 6.000 11.600 6.800 11.700 ;
        RECT 2.400 10.800 3.600 11.600 ;
        RECT 3.000 10.200 3.600 10.800 ;
        RECT 3.000 9.600 5.200 10.200 ;
        RECT 4.400 2.200 5.200 9.600 ;
        RECT 7.600 2.200 8.400 19.800 ;
        RECT 9.200 17.800 10.000 20.400 ;
        RECT 10.800 17.600 11.600 19.800 ;
        RECT 12.400 17.800 13.200 20.400 ;
        RECT 18.800 17.800 19.600 20.400 ;
        RECT 9.200 15.600 10.000 17.200 ;
        RECT 11.000 14.400 11.600 17.600 ;
        RECT 15.600 16.300 16.400 16.400 ;
        RECT 20.400 16.300 21.200 19.800 ;
        RECT 15.600 15.700 21.200 16.300 ;
        RECT 15.600 15.600 16.400 15.700 ;
        RECT 10.800 13.600 11.600 14.400 ;
        RECT 11.000 10.200 11.600 13.600 ;
        RECT 20.200 15.200 21.200 15.700 ;
        RECT 12.400 12.300 13.200 12.400 ;
        RECT 18.800 12.300 19.600 12.400 ;
        RECT 12.400 11.700 19.600 12.300 ;
        RECT 12.400 10.800 13.200 11.700 ;
        RECT 18.800 11.600 19.600 11.700 ;
        RECT 20.200 10.800 21.000 15.200 ;
        RECT 22.000 14.600 22.800 19.800 ;
        RECT 25.200 15.800 26.000 20.400 ;
        RECT 28.400 16.600 29.200 19.800 ;
        RECT 30.000 17.000 30.800 19.800 ;
        RECT 31.600 17.000 32.400 19.800 ;
        RECT 33.200 17.000 34.000 19.800 ;
        RECT 34.800 17.000 35.600 19.800 ;
        RECT 36.400 17.800 37.200 20.400 ;
        RECT 38.000 17.000 38.800 19.800 ;
        RECT 39.600 17.800 40.400 20.400 ;
        RECT 41.200 17.000 42.000 19.800 ;
        RECT 42.800 17.000 43.600 19.800 ;
        RECT 44.400 17.000 45.200 19.800 ;
        RECT 26.800 15.800 29.200 16.600 ;
        RECT 46.000 16.600 46.800 19.800 ;
        RECT 26.800 15.200 27.600 15.800 ;
        RECT 21.600 14.000 22.800 14.600 ;
        RECT 25.800 14.600 27.600 15.200 ;
        RECT 31.600 15.600 32.600 16.400 ;
        RECT 38.000 15.800 42.600 16.400 ;
        RECT 46.000 15.800 48.600 16.600 ;
        RECT 49.200 15.800 50.000 20.400 ;
        RECT 38.000 15.600 38.800 15.800 ;
        RECT 21.600 12.000 22.200 14.000 ;
        RECT 25.800 13.400 26.600 14.600 ;
        RECT 22.800 12.600 26.600 13.400 ;
        RECT 31.600 12.800 32.400 15.600 ;
        RECT 38.000 14.800 38.800 15.000 ;
        RECT 34.400 14.200 38.800 14.800 ;
        RECT 34.400 14.000 35.200 14.200 ;
        RECT 39.600 13.600 40.400 15.200 ;
        RECT 41.800 13.400 42.600 15.800 ;
        RECT 47.800 15.200 48.600 15.800 ;
        RECT 47.800 14.400 50.800 15.200 ;
        RECT 52.400 13.800 53.200 19.800 ;
        RECT 54.000 18.300 54.800 18.400 ;
        RECT 58.800 18.300 59.600 19.800 ;
        RECT 54.000 17.700 59.600 18.300 ;
        RECT 60.400 17.800 61.200 20.400 ;
        RECT 54.000 17.600 54.800 17.700 ;
        RECT 34.800 12.600 38.000 13.400 ;
        RECT 41.800 12.600 43.800 13.400 ;
        RECT 44.400 13.000 53.200 13.800 ;
        RECT 28.400 12.000 29.200 12.600 ;
        RECT 46.000 12.000 46.800 12.400 ;
        RECT 49.200 12.000 50.000 12.400 ;
        RECT 51.000 12.000 51.800 12.200 ;
        RECT 21.600 11.400 22.400 12.000 ;
        RECT 28.400 11.400 51.800 12.000 ;
        RECT 10.800 9.400 12.600 10.200 ;
        RECT 20.200 10.000 21.200 10.800 ;
        RECT 11.800 2.200 12.600 9.400 ;
        RECT 20.400 2.200 21.200 10.000 ;
        RECT 21.800 9.600 22.400 11.400 ;
        RECT 21.800 9.000 30.800 9.600 ;
        RECT 21.800 7.400 22.400 9.000 ;
        RECT 30.000 8.800 30.800 9.000 ;
        RECT 33.200 9.000 41.800 9.600 ;
        RECT 33.200 8.800 34.000 9.000 ;
        RECT 25.000 7.600 27.600 8.400 ;
        RECT 21.800 6.800 24.400 7.400 ;
        RECT 23.600 2.200 24.400 6.800 ;
        RECT 26.800 2.200 27.600 7.600 ;
        RECT 28.200 6.800 32.400 7.600 ;
        RECT 30.000 2.200 30.800 5.000 ;
        RECT 31.600 2.200 32.400 5.000 ;
        RECT 33.200 2.200 34.000 5.000 ;
        RECT 34.800 2.200 35.600 8.400 ;
        RECT 38.000 7.600 40.600 8.400 ;
        RECT 41.200 8.200 41.800 9.000 ;
        RECT 42.800 9.400 43.600 9.600 ;
        RECT 42.800 9.000 48.200 9.400 ;
        RECT 42.800 8.800 49.000 9.000 ;
        RECT 47.600 8.200 49.000 8.800 ;
        RECT 41.200 7.600 47.000 8.200 ;
        RECT 50.000 8.000 51.600 8.800 ;
        RECT 50.000 7.600 50.600 8.000 ;
        RECT 38.000 2.200 38.800 7.000 ;
        RECT 41.200 2.200 42.000 7.000 ;
        RECT 46.400 6.800 50.600 7.600 ;
        RECT 52.400 7.400 53.200 13.000 ;
        RECT 51.200 6.800 53.200 7.400 ;
        RECT 42.800 2.200 43.600 5.000 ;
        RECT 44.400 2.200 45.200 5.000 ;
        RECT 47.600 2.200 48.400 6.800 ;
        RECT 51.200 6.200 51.800 6.800 ;
        RECT 50.800 5.600 51.800 6.200 ;
        RECT 50.800 2.200 51.600 5.600 ;
        RECT 58.800 2.200 59.600 17.700 ;
      LAYER via1 ;
        RECT 6.000 25.600 6.800 26.400 ;
        RECT 34.800 34.400 35.600 35.200 ;
        RECT 38.000 35.000 38.800 35.800 ;
        RECT 33.200 32.400 34.000 33.200 ;
        RECT 23.400 29.600 24.200 30.400 ;
        RECT 20.400 23.600 21.200 24.400 ;
        RECT 42.800 27.600 43.600 28.400 ;
        RECT 33.200 24.200 34.000 25.000 ;
        RECT 34.800 24.200 35.600 25.000 ;
        RECT 36.400 24.200 37.200 25.000 ;
        RECT 38.000 24.200 38.800 25.000 ;
        RECT 41.200 24.200 42.000 25.000 ;
        RECT 44.400 24.200 45.200 25.000 ;
        RECT 46.000 24.200 46.800 25.000 ;
        RECT 47.600 24.200 48.400 25.000 ;
        RECT 7.600 13.600 8.400 14.400 ;
        RECT 38.000 14.200 38.800 15.000 ;
        RECT 49.200 11.600 50.000 12.400 ;
        RECT 31.600 6.800 32.400 7.600 ;
        RECT 34.800 6.200 35.600 7.000 ;
        RECT 30.000 4.200 30.800 5.000 ;
        RECT 31.600 4.200 32.400 5.000 ;
        RECT 33.200 4.200 34.000 5.000 ;
        RECT 38.000 6.200 38.800 7.000 ;
        RECT 41.200 6.200 42.000 7.000 ;
        RECT 42.800 4.200 43.600 5.000 ;
        RECT 44.400 4.200 45.200 5.000 ;
      LAYER metal2 ;
        RECT 6.000 29.600 6.800 30.400 ;
        RECT 9.200 29.600 10.000 30.400 ;
        RECT 17.200 29.600 18.000 30.400 ;
        RECT 23.400 29.600 24.400 30.400 ;
        RECT 6.000 27.600 6.800 28.400 ;
        RECT 15.600 27.600 16.400 28.400 ;
        RECT 6.100 26.400 6.700 27.600 ;
        RECT 6.000 25.600 6.800 26.400 ;
        RECT 9.200 25.600 10.000 26.400 ;
        RECT 6.100 16.400 6.700 25.600 ;
        RECT 9.300 16.400 9.900 25.600 ;
        RECT 10.800 19.600 11.600 20.400 ;
        RECT 10.900 18.400 11.500 19.600 ;
        RECT 10.800 17.600 11.600 18.400 ;
        RECT 15.700 16.400 16.300 27.600 ;
        RECT 20.400 23.600 21.200 24.400 ;
        RECT 33.200 24.200 34.000 37.800 ;
        RECT 34.800 24.200 35.600 37.800 ;
        RECT 36.400 24.200 37.200 37.800 ;
        RECT 38.000 24.200 38.800 35.800 ;
        RECT 41.200 24.200 42.000 35.800 ;
        RECT 42.800 27.600 43.600 28.400 ;
        RECT 6.000 15.600 6.800 16.400 ;
        RECT 9.200 15.600 10.000 16.400 ;
        RECT 15.600 15.600 16.400 16.400 ;
        RECT 6.100 12.400 6.700 15.600 ;
        RECT 7.600 13.600 8.400 14.400 ;
        RECT 6.000 11.600 6.800 12.400 ;
        RECT 18.800 12.300 19.600 12.400 ;
        RECT 20.500 12.300 21.100 23.600 ;
        RECT 42.900 20.400 43.500 27.600 ;
        RECT 44.400 24.200 45.200 35.800 ;
        RECT 46.000 24.200 46.800 37.800 ;
        RECT 47.600 24.200 48.400 37.800 ;
        RECT 49.200 29.600 50.000 30.400 ;
        RECT 54.000 29.600 54.800 30.400 ;
        RECT 42.800 19.600 43.600 20.400 ;
        RECT 18.800 11.700 21.100 12.300 ;
        RECT 18.800 11.600 19.600 11.700 ;
        RECT 30.000 4.200 30.800 17.800 ;
        RECT 31.600 4.200 32.400 17.800 ;
        RECT 33.200 4.200 34.000 17.800 ;
        RECT 34.800 6.200 35.600 17.800 ;
        RECT 38.000 6.200 38.800 17.800 ;
        RECT 39.600 13.600 40.400 14.400 ;
        RECT 41.200 6.200 42.000 17.800 ;
        RECT 42.800 4.200 43.600 17.800 ;
        RECT 44.400 4.200 45.200 17.800 ;
        RECT 49.300 12.400 49.900 29.600 ;
        RECT 54.100 18.400 54.700 29.600 ;
        RECT 54.000 17.600 54.800 18.400 ;
        RECT 49.200 11.600 50.000 12.400 ;
      LAYER via2 ;
        RECT 23.600 29.600 24.400 30.400 ;
      LAYER metal3 ;
        RECT 6.000 30.300 6.800 30.400 ;
        RECT 9.200 30.300 10.000 30.400 ;
        RECT 17.200 30.300 18.000 30.400 ;
        RECT 23.600 30.300 24.400 30.400 ;
        RECT 6.000 29.700 24.400 30.300 ;
        RECT 6.000 29.600 6.800 29.700 ;
        RECT 9.200 29.600 10.000 29.700 ;
        RECT 17.200 29.600 18.000 29.700 ;
        RECT 23.600 29.600 24.400 29.700 ;
        RECT 6.000 28.300 6.800 28.400 ;
        RECT 15.600 28.300 16.400 28.400 ;
        RECT 6.000 27.700 16.400 28.300 ;
        RECT 6.000 27.600 6.800 27.700 ;
        RECT 15.600 27.600 16.400 27.700 ;
        RECT 10.800 20.300 11.600 20.400 ;
        RECT 42.800 20.300 43.600 20.400 ;
        RECT 10.800 19.700 43.600 20.300 ;
        RECT 10.800 19.600 11.600 19.700 ;
        RECT 42.800 19.600 43.600 19.700 ;
        RECT 7.600 14.300 8.400 14.400 ;
        RECT 39.600 14.300 40.400 14.400 ;
        RECT 7.600 13.700 40.400 14.300 ;
        RECT 7.600 13.600 8.400 13.700 ;
        RECT 39.600 13.600 40.400 13.700 ;
  END
END counter
END LIBRARY

