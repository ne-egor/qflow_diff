* NGSPICE file created from counter.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

.subckt counter vdd clk rst val[0] val[1]
XFILL_0_0_0 INVX1_2/gnd vdd FILL
XFILL_0_0_1 INVX1_2/gnd vdd FILL
XFILL_0_0_2 INVX1_2/gnd vdd FILL
XBUFX2_1 INVX1_1/A INVX1_2/gnd val[0] vdd BUFX2
XBUFX2_2 DFFSR_2/Q INVX1_2/gnd val[1] vdd BUFX2
XNOR2X1_1 INVX1_1/A DFFSR_2/Q INVX1_2/gnd NOR2X1_2/A vdd NOR2X1
XNOR2X1_2 NOR2X1_2/A NOR2X1_2/B INVX1_2/gnd DFFSR_2/D vdd NOR2X1
XFILL_0_1_0 INVX1_2/gnd vdd FILL
XFILL_0_1_1 INVX1_2/gnd vdd FILL
XFILL_0_1_2 INVX1_2/gnd vdd FILL
XFILL_1_0_0 INVX1_2/gnd vdd FILL
XFILL_1_0_1 INVX1_2/gnd vdd FILL
XFILL_1_0_2 INVX1_2/gnd vdd FILL
XDFFSR_1 INVX1_1/A clk INVX1_2/Y vdd INVX1_1/Y INVX1_2/gnd vdd DFFSR
XDFFSR_2 DFFSR_2/Q clk INVX1_2/Y vdd DFFSR_2/D INVX1_2/gnd vdd DFFSR
XAND2X2_1 INVX1_1/A DFFSR_2/Q INVX1_2/gnd NOR2X1_2/B vdd AND2X2
XINVX1_1 INVX1_1/A INVX1_2/gnd INVX1_1/Y vdd INVX1
XINVX1_2 rst INVX1_2/gnd INVX1_2/Y vdd INVX1
.ends

